library verilog;
use verilog.vl_types.all;
entity Prac7_vlg_vec_tst is
end Prac7_vlg_vec_tst;
